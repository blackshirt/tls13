module tls13

fn test_extensionlist_pack_unpack_from_serverhello() ! {
	data := [u8(0x00), 0x2e, 0x00, 0x2b, 0x00, 0x02, 0x03, 0x04, 0x00, 0x33, 0x00, 0x24, 0x00,
		0x1d, 0x00, 0x20, 0x9f, 0xd7, 0xad, 0x6d, 0xcf, 0xf4, 0x29, 0x8d, 0xd3, 0xf9, 0x6d, 0x5b,
		0x1b, 0x2a, 0xf9, 0x10, 0xa0, 0x53, 0x5b, 0x14, 0x88, 0xd7, 0xf8, 0xfa, 0xbb, 0x34, 0x9a,
		0x98, 0x28, 0x80, 0xb6, 0x15]

	exts := ExtensionList.unpack(data)!
	assert exts.len == 2
	assert exts[0].tipe == .supported_versions
	ver := ProtoVersion.unpack(exts[0].data)!
	assert ver == tls_v13

	assert exts[1].tipe == .key_share
	ksh := KeyShareExtension.unpack_from_extension(exts[1], .server_hello, false)!
	assert ksh.server_share.group == .x25519
	assert ksh.server_share.key_exchange.len == 32
}
