module tls13

fn test_servernameextension_pack_unpack() ! {
	data := [u8(0x00), 0x00, 0x00, 0x18, 0x00, 0x16, 0x00, 0x00, 0x13, 0x65, 0x78, 0x61, 0x6d,
		0x70, 0x6c, 0x65, 0x2e, 0x75, 0x6c, 0x66, 0x68, 0x65, 0x69, 0x6d, 0x2e, 0x6e, 0x65, 0x74]

	sn_ext := ServerNameList.unpack_from_extension(data)!
	assert sn_ext.len == 1
	assert sn_ext[0].name_type == .host_name
	assert sn_ext[0].name.len == 0x13 // 19
	assert sn_ext[0].name.bytestr() == 'example.ulfheim.net'
}
