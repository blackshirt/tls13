module tls13

fn test_keyshareclienthello_pack_unpack() ! {
	data := [u8(0x00), 0x24, 0x00, 0x1d, 0x00, 0x20, 0x35, 0x80, 0x72, 0xd6, 0x36, 0x58, 0x80,
		0xd1, 0xae, 0xea, 0x32, 0x9a, 0xdf, 0x91, 0x21, 0x38, 0x38, 0x51, 0xed, 0x21, 0xa2, 0x8e,
		0x3b, 0x75, 0xe9, 0x65, 0xd0, 0xd2, 0xcd, 0x16, 0x62, 0x54]
	ksch := KeyShareExtension.unpack_from_extension_payload(data, .client_hello, false)!
	assert ksch.client_shares.len == 1

	ng1 := ksch.client_shares[0]
	assert ng1.group == .x25519
	assert ng1.key_exchange.len == 32

	back := ksch.pack()!
	assert back == data
}

fn test_keyshareextension_pack_unpack_for_clienthello() ! {
	data := [u8(0x00), 0x33, 0x00, 0x26, 0x00, 0x24, 0x00, 0x1d, 0x00, 0x20, 0x35, 0x80, 0x72,
		0xd6, 0x36, 0x58, 0x80, 0xd1, 0xae, 0xea, 0x32, 0x9a, 0xdf, 0x91, 0x21, 0x38, 0x38, 0x51,
		0xed, 0x21, 0xa2, 0x8e, 0x3b, 0x75, 0xe9, 0x65, 0xd0, 0xd2, 0xcd, 0x16, 0x62, 0x54]
	// test with raw extension
	ext := Extension.unpack(data)!
	assert ext.tipe == .key_share
	assert ext.length == 38
	assert ext.data.len == 38

	// test with KeyShareExtension
	out := KeyShareExtension.unpack(data, .client_hello, false)!
	assert out.msg_type == .client_hello
	assert out.is_hrr == false

	// see https://tls13.xargs.org/#client-hello/annotated
	assert out.client_shares.len == 1
	assert out.client_shares[0].group == .x25519
	assert out.client_shares[0].key_exchange == [u8(0x35), 0x80, 0x72, 0xd6, 0x36, 0x58, 0x80,
		0xd1, 0xae, 0xea, 0x32, 0x9a, 0xdf, 0x91, 0x21, 0x38, 0x38, 0x51, 0xed, 0x21, 0xa2, 0x8e,
		0x3b, 0x75, 0xe9, 0x65, 0xd0, 0xd2, 0xcd, 0x16, 0x62, 0x54]

	// pack back
	ks_ext := out.pack_to_extension()!
	back := ks_ext.pack()!
	assert back == data
}

// https://tls13.xargs.org/#server-hello
fn test_keyshareextension_pack_unpack_for_serverhello() ! {
	data := [u8(0x00), 0x33, 0x00, 0x24, 0x00, 0x1d, 0x00, 0x20, 0x9f, 0xd7, 0xad, 0x6d, 0xcf,
		0xf4, 0x29, 0x8d, 0xd3, 0xf9, 0x6d, 0x5b, 0x1b, 0x2a, 0xf9, 0x10, 0xa0, 0x53, 0x5b, 0x14,
		0x88, 0xd7, 0xf8, 0xfa, 0xbb, 0x34, 0x9a, 0x98, 0x28, 0x80, 0xb6, 0x15]

	// test with KeyShareExtension
	out := KeyShareExtension.unpack(data, .server_hello, false)!
	assert out.msg_type == .server_hello
	assert out.is_hrr == false

	assert out.server_share.group == .x25519
	assert out.server_share.key_exchange == [u8(0x9f), 0xd7, 0xad, 0x6d, 0xcf, 0xf4, 0x29, 0x8d,
		0xd3, 0xf9, 0x6d, 0x5b, 0x1b, 0x2a, 0xf9, 0x10, 0xa0, 0x53, 0x5b, 0x14, 0x88, 0xd7, 0xf8,
		0xfa, 0xbb, 0x34, 0x9a, 0x98, 0x28, 0x80, 0xb6, 0x15]

	// pack back
	back := out.pack_to_extension_bytes()!
	assert back == data
}
