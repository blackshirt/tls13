module tls13

const max_u24 = 1 << 24 - 1
