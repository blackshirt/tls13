module tls13

import encoding.binary
import crypto.rand
import blackshirt.ecdhe

// rfc 8448
const client_finished_record = [u8(0x17), 0x03, 0x03, 0x00, 0x35, 0x75, 0xec, 0x4d, 0xc2, 0x38,
	0xcc, 0xe6, 0x0b, 0x29, 0x80, 0x44, 0xa7, 0x1e, 0x21, 0x9c, 0x56, 0xcc, 0x77, 0xb0, 0x51, 0x7f,
	0xe9, 0xb9, 0x3c, 0x7a, 0x4b, 0xfc, 0x44, 0xd8, 0x7f, 0x38, 0xf8, 0x03, 0x38, 0xac, 0x98, 0xfc,
	0x46, 0xde, 0xb3, 0x84, 0xbd, 0x1c, 0xae, 0xac, 0xab, 0x68, 0x67, 0xd7, 0x26, 0xc4, 0x05, 0x46]

fn test_unpack_tls13_finished_record() ! {
	rec := TLSRecord.unpack(tls13.client_finished_record)!
	assert rec.length == 53
	assert rec.ctn_type == .application_data
}

fn test_from_openssl_output_read() ! {
	data := [u8(0x16), 0x03, 0x03, 0x00, 0x8c, 0x03, 0x03, 0x70, 0x21, 0xb1, 0x3a, 0xd7, 0x68,
		0xe7, 0x03, 0x62, 0x3a, 0xa7, 0xb5, 0x25, 0x04, 0x6f, 0xd1, 0xba, 0x83, 0x8c, 0x3e, 0xbd,
		0x73, 0xa9, 0x47, 0xed, 0x1a, 0x5c, 0x03, 0x4e, 0x09, 0x0b, 0xaa, 0x20, 0xd2, 0xfe, 0x20,
		0x1c, 0xc8, 0xe6, 0x52, 0xd8, 0x47, 0x43, 0xbf, 0xf0, 0x32, 0x6c, 0x21, 0x2f, 0x0e, 0x4d,
		0x33, 0xa3, 0xc4, 0x31, 0x25, 0xd4, 0x79, 0x34, 0x48, 0x9e, 0xef, 0x8c, 0xd8, 0x90, 0x00,
		0x02, 0x13, 0x03, 0x01, 0x00, 0x00, 0x41, 0x00, 0x0d, 0x00, 0x04, 0x00, 0x02, 0x08, 0x07,
		0x00, 0x2b, 0x00, 0x03, 0x02, 0x03, 0x04, 0x00, 0x0a, 0x00, 0x04, 0x00, 0x02, 0x00, 0x1d,
		0x00, 0x33, 0x00, 0x26, 0x00, 0x24, 0x00, 0x1d, 0x00, 0x20, 0x68, 0x04, 0xbb, 0xf7, 0xf5,
		0xa9, 0x61, 0xc4, 0xa8, 0xa1, 0x99, 0x8b, 0x68, 0x56, 0xe3, 0xd1, 0xad, 0x04, 0xa3, 0xa7,
		0x91, 0x5b, 0x1b, 0xe9, 0x94, 0x2a, 0x94, 0x88, 0xcf, 0x55, 0x83, 0x39]
	rec := TLSRecord.unpack(data)!
	// dump(rec)
}

fn test_session_init() ! {
	mut exchanger := ecdhe.new_exchanger(ecdhe.Curve.x25519)!
	// build needed random bytes
	privkey := exchanger.generate_private_key()!
	pubkey := exchanger.public_key(privkey)!

	random := rand.read(32)!
	sessid := []u8{}
	ciphersuites := [CipherSuite.tls_chacha20_poly1305_sha256]

	mut exts := []Extension{}
	// server_name extension
	srvname := new_server_name('localhost')!
	srvname_list := ServerNameList([srvname])
	srvname_ext := srvname_list.pack_to_extension()!
	exts.append(srvname_ext)

	// SupportedVersions extension
	spv := ClientSpV{
		versions: [tls_v13]
	}
	spv_ext := SupportedVersions(spv).pack_to_extension()!
	exts.append(spv_ext)

	// NamedGroupList
	ngl := NamedGroupList([NamedGroup.x25519])
	ngl_ext := ngl.pack_to_extension()!
	exts.append(ngl_ext)

	// signaturescheme
	signs_list := SignatureSchemeList([SignatureScheme.ed25519])
	signs_ext := signs_list.pack_to_extension()!
	exts.append(signs_ext)

	// KeyShare extension
	ke_entry0 := KeyShareEntry{
		group: .x25519
		key_exchange: pubkey.bytes()!
	}

	ks := KeyShareExtension{
		msg_type: .client_hello
		is_hrr: false
		client_shares: [ke_entry0]
	}
	ks_ext := ks.pack_to_extension()!
	exts.append(ks_ext)
	// TODO: add another supported extension
	ch := ClientHello{
		random: random
		legacy_session_id: sessid
		cipher_suites: ciphersuites
		extensions: exts
	}

	hsk := HandshakePayload(ch).pack_to_handshake()!
	// dump(hsk)
	pxt := TLSPlaintext.from_handshake(hsk)!
	// dump(pxt)

	pxt_obj := pxt.pack()!

	pxt_unpacked := TLSPlaintext.unpack(pxt_obj)!
	assert pxt == pxt_unpacked
	assert pxt_unpacked.ctn_type == .handshake
	assert pxt_unpacked.legacy_version == tls_v12

	hsk_unpacked := Handshake.unpack(pxt_unpacked.fragment)!
	assert hsk_unpacked.msg_type == .client_hello

	ch_unpacked := ClientHello.unpack(hsk_unpacked.payload)!
	assert ch_unpacked == ch
}

fn test_decrypted_data_from_handshake() {
	encrypted_record := [u8(233), 85, 239, 170, 3, 176, 70, 17, 90, 239, 247, 248, 245, 63, 222,
		40, 138, 128, 207, 31, 251, 196, 51]
	client_hwkey := [u8(238), 106, 116, 243, 11, 38, 234, 25, 255, 244, 246, 236, 67, 226, 151,
		139, 138, 236, 51, 254, 245, 119, 202, 186, 55, 204, 254, 223, 163, 149, 42, 244]
	client_hwiv := [u8(103), 160, 169, 56, 160, 230, 106, 13, 105, 82, 149, 5]
	server_hwkey := [u8(234), 164, 3, 81, 193, 130, 74, 52, 237, 133, 44, 180, 69, 28, 41, 81,
		18, 193, 7, 199, 68, 88, 66, 114, 106, 44, 165, 124, 126, 60, 148, 167]
	server_hwiv := [u8(24), 147, 74, 228, 50, 185, 46, 107, 41, 28, 17, 64]

	cxt := TLSCiphertext{
		opaque_type: .application_data
		legacy_version: tls_v12
		length: 23
		encrypted_record: encrypted_record
	}
	mut rc := new_record_layer(.tls_chacha20_poly1305_sha256)!
	snonce := rc.build_read_nonce(server_hwiv)
	cnonce := rc.build_read_nonce(client_hwiv)

	mut add := cxt.opaque_type.pack()!
	add << cxt.legacy_version.pack()!
	mut length := []u8{len: 2}
	binary.big_endian_put_u16(mut length, u16(cxt.length))
	add << length
	cxt_len := cxt.encrypted_record.len
	ciphertext := cxt.encrypted_record[0..cxt_len - rc.cipher.tag_size()].clone()
	plain, tag := rc.cipher.decrypt(server_hwkey, cnonce, add, ciphertext)!

	innertext := TLSInnerPlaintext.unpack(plain)!
	pxt := innertext.to_plaintext()!

	// TODO: need fix
	// dump(pxt)
}

fn test_find_content_type_position() {
	data := [u8(0), 8, 117, 139, 70, 22, 0, 0, 0, 0]
	pos := find_content_type_position(data)!
	assert pos == 5
	out := TLSInnerPlaintext.unpack(data)!
	assert out.ctn_type == .handshake
}

fn test_ee_encrypt_decrypt() {
	ee_data := [u8(0x08), 0x00, 0x00, 0x02, 0x00, 0x00]
	hsk := Handshake.unpack(ee_data)!
	assert hsk.msg_type == .encrypted_extensions
	assert hsk.length == 2
	ee := EncryptedExtensions.unpack(hsk.payload)!
	assert ee.extensions.len == 0

	client_hwkey := [u8(238), 106, 116, 243, 11, 38, 234, 25, 255, 244, 246, 236, 67, 226, 151,
		139, 138, 236, 51, 254, 245, 119, 202, 186, 55, 204, 254, 223, 163, 149, 42, 244]
	client_hwiv := [u8(103), 160, 169, 56, 160, 230, 106, 13, 105, 82, 149, 5]
	server_hwkey := [u8(234), 164, 3, 81, 193, 130, 74, 52, 237, 133, 44, 180, 69, 28, 41, 81,
		18, 193, 7, 199, 68, 88, 66, 114, 106, 44, 165, 124, 126, 60, 148, 167]
	server_hwiv := [u8(24), 147, 74, 228, 50, 185, 46, 107, 41, 28, 17, 64]

	mut rc := new_record_layer(.tls_chacha20_poly1305_sha256)!
	snonce := rc.build_read_nonce(server_hwiv)
	cnonce := rc.build_read_nonce(client_hwiv)

	pxt := TLSPlaintext.from_handshake(hsk)!
	inner := pxt.to_innerplaintext_with_padmode(.nopad)!
	plaintext := inner.pack()!
	assert plaintext.len == 7
	length := plaintext.len + rc.cipher.tag_size()

	add := rc.make_additional_data(ContentType.application_data, tls_v12, length)!
	ciphertext, tag := rc.cipher.encrypt(server_hwkey, snonce, add, plaintext)!

	mut encrypted_record := []u8{}
	encrypted_record << ciphertext
	encrypted_record << tag
	trec := TLSCiphertext{
		opaque_type: .application_data
		legacy_version: tls_v12
		length: 23
		encrypted_record: encrypted_record
	}

	txrec := rc.encrypt(pxt, server_hwkey, snonce)!
	assert trec == txrec
	cxt := trec.encrypted_record[0..trec.encrypted_record.len - rc.cipher.tag_size()]
	assert cxt == ciphertext
	dcc, mcc := rc.cipher.decrypt(server_hwkey, snonce, add, cxt)!
	dec_trec := rc.decrypt(trec, server_hwkey, server_hwiv)!

	assert dcc == plaintext
	assert dec_trec == pxt
	assert tag == mcc

	dcc_inn := TLSInnerPlaintext.unpack(dcc)!
	exx := dcc_inn.to_plaintext()!

	eex := Handshake.unpack(exx.fragment)!
	assert eex.msg_type == .encrypted_extensions
	assert eex.length == 2
}

fn test_certificate_msg_from_session() ! {
	cert_msg := [u8(0x0b), 0x00, 0x01, 0xac, 0x00, 0x00, 0x01, 0xa8, 0x00, 0x01, 0xa3, 0x30, 0x82,
		0x01, 0x9f, 0x30, 0x82, 0x01, 0x51, 0xa0, 0x03, 0x02, 0x01, 0x02, 0x02, 0x14, 0x7f, 0xe5,
		0x3c, 0xfb, 0x10, 0x10, 0x61, 0x40, 0xd3, 0xe7, 0xde, 0xfb, 0xe3, 0x4f, 0xc0, 0xfa, 0x20,
		0xcc, 0xa8, 0x03, 0x30, 0x05, 0x06, 0x03, 0x2b, 0x65, 0x70, 0x30, 0x45, 0x31, 0x0b, 0x30,
		0x09, 0x06, 0x03, 0x55, 0x04, 0x06, 0x13, 0x02, 0x41, 0x55, 0x31, 0x13, 0x30, 0x11, 0x06,
		0x03, 0x55, 0x04, 0x08, 0x0c, 0x0a, 0x53, 0x6f, 0x6d, 0x65, 0x2d, 0x53, 0x74, 0x61, 0x74,
		0x65, 0x31, 0x21, 0x30, 0x1f, 0x06, 0x03, 0x55, 0x04, 0x0a, 0x0c, 0x18, 0x49, 0x6e, 0x74,
		0x65, 0x72, 0x6e, 0x65, 0x74, 0x20, 0x57, 0x69, 0x64, 0x67, 0x69, 0x74, 0x73, 0x20, 0x50,
		0x74, 0x79, 0x20, 0x4c, 0x74, 0x64, 0x30, 0x1e, 0x17, 0x0d, 0x32, 0x33, 0x31, 0x31, 0x31,
		0x33, 0x31, 0x33, 0x32, 0x30, 0x30, 0x39, 0x5a, 0x17, 0x0d, 0x32, 0x34, 0x31, 0x31, 0x31,
		0x32, 0x31, 0x33, 0x32, 0x30, 0x30, 0x39, 0x5a, 0x30, 0x45, 0x31, 0x0b, 0x30, 0x09, 0x06,
		0x03, 0x55, 0x04, 0x06, 0x13, 0x02, 0x41, 0x55, 0x31, 0x13, 0x30, 0x11, 0x06, 0x03, 0x55,
		0x04, 0x08, 0x0c, 0x0a, 0x53, 0x6f, 0x6d, 0x65, 0x2d, 0x53, 0x74, 0x61, 0x74, 0x65, 0x31,
		0x21, 0x30, 0x1f, 0x06, 0x03, 0x55, 0x04, 0x0a, 0x0c, 0x18, 0x49, 0x6e, 0x74, 0x65, 0x72,
		0x6e, 0x65, 0x74, 0x20, 0x57, 0x69, 0x64, 0x67, 0x69, 0x74, 0x73, 0x20, 0x50, 0x74, 0x79,
		0x20, 0x4c, 0x74, 0x64, 0x30, 0x2a, 0x30, 0x05, 0x06, 0x03, 0x2b, 0x65, 0x70, 0x03, 0x21,
		0x00, 0xbd, 0xe2, 0xcf, 0x61, 0x4b, 0xa2, 0x71, 0x81, 0x67, 0x06, 0x21, 0x9a, 0x26, 0xc5,
		0x94, 0x3f, 0x1c, 0x98, 0x2d, 0x93, 0x33, 0x0a, 0x5b, 0x82, 0x54, 0x81, 0x3f, 0x85, 0x4f,
		0xf2, 0xdb, 0xcd, 0xa3, 0x53, 0x30, 0x51, 0x30, 0x1d, 0x06, 0x03, 0x55, 0x1d, 0x0e, 0x04,
		0x16, 0x04, 0x14, 0xdb, 0x33, 0x49, 0xb5, 0x72, 0xa3, 0x0d, 0xbc, 0xd3, 0x7d, 0x15, 0xcf,
		0xe0, 0xfb, 0xe6, 0xaa, 0xf1, 0x38, 0x05, 0xb5, 0x30, 0x1f, 0x06, 0x03, 0x55, 0x1d, 0x23,
		0x04, 0x18, 0x30, 0x16, 0x80, 0x14, 0xdb, 0x33, 0x49, 0xb5, 0x72, 0xa3, 0x0d, 0xbc, 0xd3,
		0x7d, 0x15, 0xcf, 0xe0, 0xfb, 0xe6, 0xaa, 0xf1, 0x38, 0x05, 0xb5, 0x30, 0x0f, 0x06, 0x03,
		0x55, 0x1d, 0x13, 0x01, 0x01, 0xff, 0x04, 0x05, 0x30, 0x03, 0x01, 0x01, 0xff, 0x30, 0x05,
		0x06, 0x03, 0x2b, 0x65, 0x70, 0x03, 0x41, 0x00, 0xa7, 0x45, 0xce, 0x36, 0xef, 0x28, 0x9d,
		0x81, 0xdc, 0xd1, 0x22, 0x20, 0x80, 0x25, 0xc6, 0xf2, 0x50, 0x53, 0xba, 0xe4, 0x98, 0x6d,
		0x04, 0xe3, 0xb4, 0xcc, 0xb6, 0x48, 0x20, 0x3f, 0x8b, 0xc8, 0x30, 0x5d, 0xed, 0x91, 0xa4,
		0xd6, 0x15, 0xc8, 0xd9, 0x6b, 0x7c, 0xb6, 0x19, 0x9b, 0x6b, 0x4d, 0xdc, 0xa5, 0x19, 0xfb,
		0xef, 0x2e, 0x50, 0x1e, 0x2b, 0xb7, 0x4c, 0x12, 0xcd, 0x41, 0x00, 0x07, 0x00, 0x00]

	cert := Handshake.unpack(cert_msg)!
	certback := cert.pack()!
	assert certback.len == 0x01b0 // 132

	assert cert_msg == certback
}
