module tls13

import encoding.binary
