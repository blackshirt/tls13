module tls13

fn test_signatureschemeextension_pack_unpack() ! {
	bytes := [u8(0x00), 0x0d, 0x00, 0x1e, 0x00, 0x1c, 0x04, 0x03, 0x05, 0x03, 0x06, 0x03, 0x08,
		0x07, 0x08, 0x08, 0x08, 0x09, 0x08, 0x0a, 0x08, 0x0b, 0x08, 0x04, 0x08, 0x05, 0x08, 0x06,
		0x04, 0x01, 0x05, 0x01, 0x06, 0x01]

	ext := Extension.unpack(bytes)!
	assert ext.tipe == .signature_algorithms
	assert ext.length == 30

	signs := SignatureSchemeList.unpack_from_extension_bytes(bytes)!
	assert signs.len == 14

	// pack back
	back := signs.pack_to_extension_bytes()!
	assert back == bytes
}
